// hex_led.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module hex_led (
		input  wire       clk_clk,                              //                            clk.clk
		input  wire [7:0] eightbitstosevenseg_0_data_in_export, //  eightbitstosevenseg_0_data_in.export
		output wire [6:0] eightbitstosevenseg_0_led_pins_led0,  // eightbitstosevenseg_0_led_pins.led0
		output wire [6:0] eightbitstosevenseg_0_led_pins_led1,  //                               .led1
		input  wire [7:0] eightbitstosevenseg_1_data_in_export, //  eightbitstosevenseg_1_data_in.export
		output wire [6:0] eightbitstosevenseg_1_led_pins_led0,  // eightbitstosevenseg_1_led_pins.led0
		output wire [6:0] eightbitstosevenseg_1_led_pins_led1,  //                               .led1
		input  wire [7:0] eightbitstosevenseg_2_data_in_export, //  eightbitstosevenseg_2_data_in.export
		output wire [6:0] eightbitstosevenseg_2_led_pins_led0,  // eightbitstosevenseg_2_led_pins.led0
		output wire [6:0] eightbitstosevenseg_2_led_pins_led1,  //                               .led1
		input  wire       reset_reset_n                         //                          reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [EightBitsToSevenSeg_0:reset, EightBitsToSevenSeg_1:reset, EightBitsToSevenSeg_2:reset]

	EightBitsToSevenSeg eightbitstosevenseg_0 (
		.hexval (eightbitstosevenseg_0_data_in_export), //  data_in.export
		.digit0 (eightbitstosevenseg_0_led_pins_led0),  // led_pins.led0
		.digit1 (eightbitstosevenseg_0_led_pins_led1),  //         .led1
		.reset  (rst_controller_reset_out_reset),       //    reset.reset
		.clock  (clk_clk)                               //    clock.clk
	);

	EightBitsToSevenSeg eightbitstosevenseg_1 (
		.hexval (eightbitstosevenseg_1_data_in_export), //  data_in.export
		.digit0 (eightbitstosevenseg_1_led_pins_led0),  // led_pins.led0
		.digit1 (eightbitstosevenseg_1_led_pins_led1),  //         .led1
		.reset  (rst_controller_reset_out_reset),       //    reset.reset
		.clock  (clk_clk)                               //    clock.clk
	);

	EightBitsToSevenSeg eightbitstosevenseg_2 (
		.hexval (eightbitstosevenseg_2_data_in_export), //  data_in.export
		.digit0 (eightbitstosevenseg_2_led_pins_led0),  // led_pins.led0
		.digit1 (eightbitstosevenseg_2_led_pins_led1),  //         .led1
		.reset  (rst_controller_reset_out_reset),       //    reset.reset
		.clock  (clk_clk)                               //    clock.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
